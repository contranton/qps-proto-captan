package ads9813_pkg is

subtype t_ADS9813_DATA_RATE is integer range 1 to 2;

end package ads9813_pkg;

package body ads9813_pkg is


end package body ads9813_pkg;
