library ieee;
use ieee.numeric_std.all;

package sim_pkg is

 subtype t_FREQUENCY_MHZ is real;

end package sim_pkg;
